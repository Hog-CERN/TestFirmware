LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY example;
LIBRARY xil_defaultlib;
USE xil_defaultlib.all;

ENTITY TB_example_xsim IS
END TB_example_xsim;

ARCHITECTURE behavior OF TB_example_xsim IS 
    constant DATA_WIDTH : integer := 16;
    
    
    --Inputs
    signal CLK      : std_logic := '0';
    signal RST      : std_logic := '0';
    signal DataIn   : std_logic_vector(DATA_WIDTH-1 downto 0) := (others => '0');
    signal ReadEn   : std_logic := '0';
    signal WriteEn  : std_logic := '0';
    
    --Outputs
    signal DataOut  : std_logic_vector(DATA_WIDTH-1 downto 0);
    signal Empty    : std_logic;
    signal Full     : std_logic;
    
    -- Clock period definitions
    constant CLK_period : time := 10 ns;

BEGIN

    -- Instantiate the Unit Under Test (UUT)
    uut: entity xil_defaultlib.top_example
        PORT MAP (
            CLK     => CLK,
            RST     => RST,
            DataIn  => DataIn,
            WriteEn => WriteEn,
            ReadEn  => ReadEn,
            DataOut => DataOut,
            Full    => Full,
            Empty   => Empty
        );
    
    -- Clock process definitions
    CLK_process :process
    begin
        CLK <= '0';
        wait for CLK_period/2;
        CLK <= '1';
        wait for CLK_period/2;
    end process;
    
    -- Reset process
    rst_proc : process
    begin
    wait for CLK_period * 5;
        
        RST <= '1';
        
        wait for CLK_period * 5;
        
        RST <= '0';
        
        wait;
    end process;
    
    -- Write process
    wr_proc : process
        variable counter : unsigned (DATA_WIDTH-1 downto 0) := (others => '0');
    begin       
        wait for CLK_period * 20;

        for i in 1 to 32 loop
            counter := counter + 1;
            
            DataIn <= std_logic_vector(counter);
            
            wait for CLK_period * 1;
            
            WriteEn <= '1';
            
            wait for CLK_period * 1;
        
            WriteEn <= '0';
        end loop;
        
        wait for clk_period * 20;
        
        for i in 1 to 32 loop
            counter := counter + 1;
            
            DataIn <= std_logic_vector(counter);
            
            wait for CLK_period * 1;
            
            WriteEn <= '1';
            
            wait for CLK_period * 1;
            
            WriteEn <= '0';
        end loop;
        
        wait;
    end process;
    
    -- Read process
    rd_proc : process
    begin
        wait for CLK_period * 20;
        
        wait for CLK_period * 40;
            
        ReadEn <= '1';
        
        wait for CLK_period * 60;
        
        ReadEn <= '0';
        
        wait for CLK_period * 256 * 2;
        
        ReadEn <= '1';
        
        wait;
    end process;

END;
